library verilog;
use verilog.vl_types.all;
entity FPU_32b_vlg_vec_tst is
end FPU_32b_vlg_vec_tst;
