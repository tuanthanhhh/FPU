library verilog;
use verilog.vl_types.all;
entity tb_FPU_32b is
end tb_FPU_32b;
