library verilog;
use verilog.vl_types.all;
entity tb_Adder_32bit is
end tb_Adder_32bit;
